module backwards_pass
(
    // ask about how many weight abouts and shit and if i should just make hidden layer smaller to fix this 
    
)


//honestly just thug it out
//oh also i think tmrw just do lfsr method 


endmodule
