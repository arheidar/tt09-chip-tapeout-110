module hidden_backwards_pass
(
    input target_i,
    input en_i,
    //do these need to be reg?
    output hw0_o,
    output hw1_o,
    output hw2_o,
    output hw3_o,
    output hw4_o,
    output hw5_o,
    output hw6_o,
    output hw7_o,
    output ow0_o,
    output ow1_o    
);


//might just change this to be a backwards pass implemented in each neuron but idk yet


endmodule
