module hidden_backprop
(
    input target_i,
    input en_i,

    
    input [7:0] w0_i, 
    input [7:0] w1_i, 
    input [7:0] w2_i, 
    input [7:0] w3_i, 

);


//might just change this to be a backwards pass implemented in each neuron but idk yet


endmodule
