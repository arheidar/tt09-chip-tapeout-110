module state_mach
//inputs named in a x_(to)_y_i format based on my state machine diagram
    input init_f1_i,
    input f_b_i,
    input b_f2_i,
    output
    //just realized if im doing lfsr method ima need a more complex sm. ig we'll see
    


endmodule